
module SBqM;





counter counter1();
CLOCK CLK1 ; 


endmodule 